/* Verilog model created from schematic schemaSR.sch -- Mar 26, 2016 15:20 */

module schemaSR;




endmodule // schemaSR
